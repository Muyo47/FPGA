--Tu bitmap esta preparado! Copia lo siguiente:

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity ROMx2 is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(8-1 downto 0);
    dout : out std_logic_vector(16-1 downto 0));
end ROMx2;


architecture BEHAVIORAL of ROMx2 is
  signal addr_int  : natural range 0 to 2**8-1;
 type memostruct is array (natural range<>) of std_logic_vector(16-1 downto 0);
 constant filaimg : memostruct := (
 -- FONDO PLANO
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO RECTO VERTICAL
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
-- MURO RECTO HORIZONTAL
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO FIN HORIZONTAL IZQUIERDA
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000001111111111",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000001111111111",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO FIN HORIZONTAL DERECHA
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"1111111111000000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"1111111111000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO FIN VERTICAL ARRIBA
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000001111000000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
-- MURO FIN VERTICAL ABAJO
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000001111000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- GIRO ARRIBA DERECHA
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000001111111111",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000011111111000",
"0000011111110000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
-- GIRO ARRIBA IZQUIERDA
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"1111111111000000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"0001111111100000",
"0000111111100000",
"0000011111100000",
"0000011111100000",
"0000011111100000",
-- GIRO ABAJO DERECHA
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000011111110000",
"0000011111111000",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000011111111111",
"0000001111111111",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- GIRO ABAJO IZQUIERDA
"0000011111100000",
"0000011111100000",
"0000011111100000",
"0000111111100000",
"0001111111100000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"1111111111100000",
"1111111111000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- LUIGI
"0000000000000000",
"0000000000000000",
"0000011111000000",
"0000111111111000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000111111110000",
"0001111111111000",
"0011111111111100",
"0000110110110000",
"0000011111100000",
"0000111111110000",
"0000111111110000");



begin

 addr_int <= TO_INTEGER(unsigned(addr));

 P_ROM: process (clk)
  begin
   if clk'event and clk='1' then
     dout <= filaimg(addr_int);
    end if;
 end process;

end BEHAVIORAL;
