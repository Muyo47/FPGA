library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_temp is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(5-1 downto 0);
    dout : out std_logic_vector(32-1 downto 0) 
  );
end ROM_temp;


architecture BEHAVIORAL of ROM_temp is
  signal addr_int  : natural range 0 to 2**5-1;
  type memostruct is array (natural range<>) of std_logic_vector(32-1 downto 0);
  constant filaimg : memostruct := (
       "00000000000000000000000000000000",
       "11100000000000000001110000111000",
       "00000011111111110000011100000000",
       "00001111111111111000011100000000",
       "00011001111111111100000000000000",
       "00111001111111111110000000000000",
       "00111001111000111111111111100000",
       "00111001111110011111111111110000",
       "00111001011110001111111111111000",
       "00111001011110000000000011111000",
       "00111000000000111000000001111100",
       "00111000000000111000000011111100",
       "00111000000000111000000011111100",
       "00111000000000111000000011111000",
       "00111001000000000000000011100000",
       "00111001110000000000000000000000",
       "00111001111000000001110000000000",
       "00011001111100000001111111100000",
       "00001001111110001111111111110000",
       "00001001111110001111111111111000",
       "00001111111110001111111011111100",
       "00001111111110001111111011111100",
       "00001111111110001111111011111100",
       "00001111000010001111111111111100",
       "00001111000011111111111111111100",
       "00001111000011111111111111111100",
       "00001111000011111111111111111000",
       "00001111000011111111111111110000",
       "00000000001111111111000000000000",
       "00000000001111111111000000000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;