-- ROM PLANO 0

-- FONDO PLANO 0000
-- MURO RECTO VERTICAL 0001  1
-- MURO RECTO HORIZONTAL 0010  2
-- MURO FIN HORIZONTAL DERECHA 0011  3
-- MURO FIN HORIZONTAL IZQUIERDA 0100  4
-- MURO FIN VERTICAL ARRIBA 0101  5
-- MURO FIN VERTICAL ABAJO 0110  6
-- FONDO PLANO 0111  7
-- GIRO ARRIBA IZQUIERDA 1000  8
-- GIRO ARRIBA DERECHA 1001  9
-- GIRO ABAJO IZQUIERDA 1010  10
-- GIRO ABAJO DERECHA 1011  11
-- FONDO PLANO 1100  12
-- FONDO PLANO 1101  13
-- FONDO PLANO 1110  14
-- LUIGI 1111  15

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity ROMx is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(8-1 downto 0);
    dout : out std_logic_vector(16-1 downto 0));
end ROMx;


architecture BEHAVIORAL of ROMx is
  signal addr_int  : natural range 0 to 2**8-1;
 type memostruct is array (natural range<>) of std_logic_vector(16-1 downto 0);
 constant filaimg : memostruct := (
 -- FONDO PLANO 0000
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO RECTO VERTICAL 0001
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
-- MURO RECTO HORIZONTAL 0010
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO FIN HORIZONTAL IZQUIERDA 0011
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000001111111111",
"0000011111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000011111111111",
"0000001111111111",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO FIN HORIZONTAL DERECHA 0100
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"1111111111000000",
"1111111111100000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111100000",
"1111111111000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- MURO FIN VERTICAL ARRIBA 0101
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000001111000000",
"0000011111100000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
-- MURO FIN VERTICAL ABAJO 0110
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000011111100000",
"0000001111000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO 0111
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- GIRO ARRIBA DERECHA 1000
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000001111111111",
"0000011111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
-- GIRO ARRIBA IZQUIERDA 1001
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"1111111111000000",
"1111111111100000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"0001111111110000",
"0000111111110000",
"0000111111110000",
"0000111111110000",
-- GIRO ABAJO DERECHA 1010
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0000111111111000",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000111111111111",
"0000011111111111",
"0000001111111111",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- GIRO ABAJO IZQUIERDA 1011
"0000111111110000",
"0000111111110000",
"0000111111110000",
"0001111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111110000",
"1111111111100000",
"1111111111000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO 1100
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO 1101
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- FONDO PLANO 1110
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
-- LUIGI 1111
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000000000000000",
"0000111110100000",
"0001111110111000",
"0001111111011100",
"0001111110001000",
"0000011111100000",
"0000001001000000",
"0000001001000000",
"0000001111000000",
"0011011111101100",
"0011111111111100",
"0011111111111100",
"0000111111110000");


begin

 addr_int <= TO_INTEGER(unsigned(addr));

 P_ROM: process (clk)
  begin
   if clk'event and clk='1' then
     dout <= filaimg(addr_int);
    end if;
 end process;

end BEHAVIORAL;
